`ifndef _IO_MAP_INCLUDED
`define _IO_MAP_INCLUDED

`define SYS_CLK_FREQ 100

`define BRIDGE_BASE 0xc0000000

`define S0_SYS_TIMER 0
`define S1_UART1     1
`define S2_LED       2
`define S3_SW        3
`define S4_XADC      4

`endif